module elevator_top (
    input clk,rst,
    input [2:0] req_floor,
    input emergency_stop,
    output [1:0] door,
    output [2:0] current_floor,
    output [7:0] requests,
    output up,down,idle,
);


    
endmodule